module and32sb(out,a,b);
input a;
input b;
output [31:0] out;

and ad01(out[0],a,b);
and ad02(out[1],a,b);
and ad03(out[2],a,b);
and ad04(out[3],a,b);
and ad05(out[4],a,b);
and ad06(out[5],a,b);
and ad07(out[6],a,b);
and ad08(out[7],a,b);
and ad09(out[8],a,b);
and ad010(out[9],a,b);
and ad011(out[10],a,b);
and ad012(out[11],a,b);
and ad013(out[12],a,b);
and ad014(out[13],a,b);
and ad015(out[14],a,b);
and ad016(out[15],a,b);
and ad017(out[16],a,b);
and ad018(out[17],a,b);
and ad019(out[18],a,b);
and ad020(out[19],a,b);
and ad021(out[20],a,b);
and ad022(out[21],a,b);
and ad023(out[22],a,b);
and ad024(out[23],a,b);
and ad025(out[24],a,b);
and ad026(out[25],a,b);
and ad027(out[26],a,b);
and ad028(out[27],a,b);
and ad029(out[28],a,b);
and ad030(out[29],a,b);
and ad031(out[30],a,b);
and ad032(out[31],a,b);

endmodule
