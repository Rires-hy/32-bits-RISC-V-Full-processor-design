module and32(out,a,b);
input [31:0] a;
input b;
output [31:0] out;

and ad01(out[0],a[0],b);
and ad02(out[1],a[1],b);
and ad03(out[2],a[2],b);
and ad04(out[3],a[3],b);
and ad05(out[4],a[4],b);
and ad06(out[5],a[5],b);
and ad07(out[6],a[6],b);
and ad08(out[7],a[7],b);
and ad09(out[8],a[8],b);
and ad010(out[9],a[9],b);
and ad011(out[10],a[10],b);
and ad012(out[11],a[11],b);
and ad013(out[12],a[12],b);
and ad014(out[13],a[13],b);
and ad015(out[14],a[14],b);
and ad016(out[15],a[15],b);
and ad017(out[16],a[16],b);
and ad018(out[17],a[17],b);
and ad019(out[18],a[18],b);
and ad020(out[19],a[19],b);
and ad021(out[20],a[20],b);
and ad022(out[21],a[21],b);
and ad023(out[22],a[22],b);
and ad024(out[23],a[23],b);
and ad025(out[24],a[24],b);
and ad026(out[25],a[25],b);
and ad027(out[26],a[26],b);
and ad028(out[27],a[27],b);
and ad029(out[28],a[28],b);
and ad030(out[29],a[29],b);
and ad031(out[30],a[30],b);
and ad032(out[31],a[31],b);

endmodule
