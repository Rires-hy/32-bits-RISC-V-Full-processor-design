module Rshift(out,a,s);
input [31:0] a;
input [4:0] s;
output [31:0] out;

wire [31:0] w0; 
wire [31:0] w1; 
wire [31:0] w2; 
wire [31:0] w3; 
wire [31:0] w4;
wire [31:0] o0; 
wire [31:0] o1; 
wire [31:0] o2; 
wire [31:0] o3; 
wire [31:0] o4; 

wire [31:0] d;
assign d[31:0] = a[31]? {32'b11111111111111111111111111111111}: {32'b00000000000000000000000000000000};

//s[0]
assign w0[31:0]={d[0],a[31:1]};
MUX2 m0(o0[31:0],w0[31:0],a[31:0],~s[0]);

//s[1]
assign w1[31:0]={d[1:0],a[31:2]};
MUX2 m1(o1[31:0],w1[31:0],o0[31:0],~s[1]);

//s[2]
assign w2[31:0]={d[3:0],a[31:4]};
MUX2 m2(o2[31:0],w2[31:0],o1[31:0],~s[2]);

//s[3]
assign w3[31:0]={d[7:0],a[31:8]};
MUX2 m3(o3[31:0],w3[31:0],o2[31:0],~s[3]);

//s[4]
assign w4[31:0]={d[15:0],a[31:16]};
MUX2 m4(out[31:0],w4[31:0],o3[31:0],~s[4]);

endmodule
