module and32(out,a,b);
input [31:0] a;
input [31:0] b;
output [31:0] out;

and ad01(out[0],a[0],b[0]);
and ad02(out[1],a[1],b[1]);
and ad03(out[2],a[2],b[2]);
and ad04(out[3],a[3],b[3]);
and ad05(out[4],a[4],b[4]);
and ad06(out[5],a[5],b[5]);
and ad07(out[6],a[6],b[6]);
and ad08(out[7],a[7],b[7]);
and ad09(out[8],a[8],b[8]);
and ad010(out[9],a[9],b[9]);
and ad011(out[10],a[10],b[10]);
and ad012(out[11],a[11],b[11]);
and ad013(out[12],a[12],b[12]);
and ad014(out[13],a[13],b[13]);
and ad015(out[14],a[14],b[14]);
and ad016(out[15],a[15],b[15]);
and ad017(out[16],a[16],b[16]);
and ad018(out[17],a[17],b[17]);
and ad019(out[18],a[18],b[18]);
and ad020(out[19],a[19],b[19]);
and ad021(out[20],a[20],b[20]);
and ad022(out[21],a[21],b[21]);
and ad023(out[22],a[22],b[22]);
and ad024(out[23],a[23],b[23]);
and ad025(out[24],a[24],b[24]);
and ad026(out[25],a[25],b[25]);
and ad027(out[26],a[26],b[26]);
and ad028(out[27],a[27],b[27]);
and ad029(out[28],a[28],b[28]);
and ad030(out[29],a[29],b[29]);
and ad031(out[30],a[30],b[30]);
and ad032(out[31],a[31],b[31]);

endmodule
